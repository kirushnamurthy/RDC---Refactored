module tb_top();
    initial begin
        $display("Hello, SystemVerilog!");
        $finish;
    end
endmodule 